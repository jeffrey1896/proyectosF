limite_inst : limite PORT MAP (
		result	 => result_sig
	);
