uno_inst : uno PORT MAP (
		result	 => result_sig
	);
