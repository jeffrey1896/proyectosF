cinco_inst : cinco PORT MAP (
		result	 => result_sig
	);
